`timescale 1ms/1ns

module numeric_code_detonator_tb ();

initial begin
    
end

endmodule