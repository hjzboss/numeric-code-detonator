////////////////////////////////////////////////////////////////////////////////
// 公司: NUDT
// 工程师: 黄俊哲
// 创建日期: 2022/11/07
// 设计名称: 数字密码引爆器
// 模块名: key_debounce_tb
// 目标器件: 未定
// 工具软件版本号: vivado
// 描述:
// 按键消抖电路的testbench
// 修订版本:
// rev1.0
// 额外注释:
// 待定
////////////////////////////////////////////////////////////////////////////////

`timescale 1ms/1ns

module key_debounce_tb ();
    // todo
endmodule