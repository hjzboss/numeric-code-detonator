`timescale 1ms/1ns

module key_debounce_tb ();
    
endmodule